--! Standard libraries
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--! User packages
use work.tf_pkg.all;
use work.memUtil_pkg.all;

entity SectorProcessorFull is
  port(
    clk        : in std_logic;
    reset      : in std_logic;
    IR_start  : in std_logic;
    IR_bx_in : in std_logic_vector(2 downto 0);
    FT_bx_out : out std_logic_vector(2 downto 0);
    FT_bx_out_vld : out std_logic;
    FT_done   : out std_logic;
    PR_bx_out : out std_logic_vector(2 downto 0);
    PR_bx_out_vld : out std_logic;
    PR_done   : out std_logic;
    ME_bx_out : out std_logic_vector(2 downto 0);
    ME_bx_out_vld : out std_logic;
    ME_done   : out std_logic;
    MC_bx_out : out std_logic_vector(2 downto 0);
    MC_bx_out_vld : out std_logic;
    MC_done   : out std_logic;
    IR_bx_out : out std_logic_vector(2 downto 0);
    IR_bx_out_vld : out std_logic;
    IR_done   : out std_logic;
    TE_bx_out : out std_logic_vector(2 downto 0);
    TE_bx_out_vld : out std_logic;
    TE_done   : out std_logic;
    VMR_bx_out : out std_logic_vector(2 downto 0);
    VMR_bx_out_vld : out std_logic;
    VMR_done   : out std_logic;
    TC_bx_out : out std_logic_vector(2 downto 0);
    TC_bx_out_vld : out std_logic;
    TC_done   : out std_logic;
    DL_39_link_AV_dout       : in t_arr_DL_39_DATA;
    DL_39_link_empty_neg     : in t_arr_DL_39_1b;
    DL_39_link_read          : out t_arr_DL_39_1b;
    IL_36_mem_A_wea        : out t_arr_IL_36_1b;
    IL_36_mem_AV_writeaddr : out t_arr_IL_36_ADDR;
    IL_36_mem_AV_din       : out t_arr_IL_36_DATA;
    AS_36_mem_A_wea        : out t_arr_AS_36_1b;
    AS_36_mem_AV_writeaddr : out t_arr_AS_36_ADDR;
    AS_36_mem_AV_din       : out t_arr_AS_36_DATA;
    VMSME_16_mem_A_wea        : out t_arr_VMSME_16_1b;
    VMSME_16_mem_AV_writeaddr : out t_arr_VMSME_16_ADDR;
    VMSME_16_mem_AV_din       : out t_arr_VMSME_16_DATA;
    VMSME_17_mem_A_wea        : out t_arr_VMSME_17_1b;
    VMSME_17_mem_AV_writeaddr : out t_arr_VMSME_17_ADDR;
    VMSME_17_mem_AV_din       : out t_arr_VMSME_17_DATA;
    VMSTE_22_mem_A_wea        : out t_arr_VMSTE_22_1b;
    VMSTE_22_mem_AV_writeaddr : out t_arr_VMSTE_22_ADDR;
    VMSTE_22_mem_AV_din       : out t_arr_VMSTE_22_DATA;
    VMSTE_16_mem_A_wea        : out t_arr_VMSTE_16_1b;
    VMSTE_16_mem_AV_writeaddr : out t_arr_VMSTE_16_ADDR;
    VMSTE_16_mem_AV_din       : out t_arr_VMSTE_16_DATA;
    SP_14_mem_A_wea        : out t_arr_SP_14_1b;
    SP_14_mem_AV_writeaddr : out t_arr_SP_14_ADDR;
    SP_14_mem_AV_din       : out t_arr_SP_14_DATA;
    TPROJ_60_mem_A_wea        : out t_arr_TPROJ_60_1b;
    TPROJ_60_mem_AV_writeaddr : out t_arr_TPROJ_60_ADDR;
    TPROJ_60_mem_AV_din       : out t_arr_TPROJ_60_DATA;
    TPROJ_58_mem_A_wea        : out t_arr_TPROJ_58_1b;
    TPROJ_58_mem_AV_writeaddr : out t_arr_TPROJ_58_ADDR;
    TPROJ_58_mem_AV_din       : out t_arr_TPROJ_58_DATA;
    TPAR_70_mem_A_wea        : out t_arr_TPAR_70_1b;
    TPAR_70_mem_AV_writeaddr : out t_arr_TPAR_70_ADDR;
    TPAR_70_mem_AV_din       : out t_arr_TPAR_70_DATA;
    VMPROJ_24_mem_A_wea        : out t_arr_VMPROJ_24_1b;
    VMPROJ_24_mem_AV_writeaddr : out t_arr_VMPROJ_24_ADDR;
    VMPROJ_24_mem_AV_din       : out t_arr_VMPROJ_24_DATA;
    AP_60_mem_A_wea        : out t_arr_AP_60_1b;
    AP_60_mem_AV_writeaddr : out t_arr_AP_60_ADDR;
    AP_60_mem_AV_din       : out t_arr_AP_60_DATA;
    AP_58_mem_A_wea        : out t_arr_AP_58_1b;
    AP_58_mem_AV_writeaddr : out t_arr_AP_58_ADDR;
    AP_58_mem_AV_din       : out t_arr_AP_58_DATA;
    CM_14_mem_A_wea        : out t_arr_CM_14_1b;
    CM_14_mem_AV_writeaddr : out t_arr_CM_14_ADDR;
    CM_14_mem_AV_din       : out t_arr_CM_14_DATA;
    FM_52_mem_A_wea        : out t_arr_FM_52_1b;
    FM_52_mem_AV_writeaddr : out t_arr_FM_52_ADDR;
    FM_52_mem_AV_din       : out t_arr_FM_52_DATA;
    TW_84_stream_AV_din       : out t_arr_TW_84_DATA;
    TW_84_stream_A_full_neg   : in t_arr_TW_84_1b;
    TW_84_stream_A_write      : out t_arr_TW_84_1b;
    BW_46_stream_AV_din       : out t_arr_BW_46_DATA;
    BW_46_stream_A_full_neg   : in t_arr_BW_46_1b;
    BW_46_stream_A_write      : out t_arr_BW_46_1b
  );
end SectorProcessorFull;

architecture rtl of SectorProcessorFull is

  signal IL_36_mem_A_enb          : t_arr_IL_36_1b;
  signal IL_36_mem_AV_readaddr    : t_arr_IL_36_ADDR;
  signal IL_36_mem_AV_dout        : t_arr_IL_36_DATA;
  signal IL_36_mem_AAV_dout_nent  : t_arr_IL_36_NENT; -- (#page)
  signal AS_36_mem_A_enb          : t_arr_AS_36_1b;
  signal AS_36_mem_AV_readaddr    : t_arr_AS_36_ADDR;
  signal AS_36_mem_AV_dout        : t_arr_AS_36_DATA;
  signal VMSME_16_mem_A_enb          : t_arr_VMSME_16_1b;
  signal VMSME_16_mem_AV_readaddr    : t_arr_VMSME_16_ADDR;
  signal VMSME_16_mem_AV_dout        : t_arr_VMSME_16_DATA;
  signal VMSME_16_mem_AAAV_dout_nent : t_arr_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_17_mem_A_enb          : t_arr_VMSME_17_1b;
  signal VMSME_17_mem_AV_readaddr    : t_arr_VMSME_17_ADDR;
  signal VMSME_17_mem_AV_dout        : t_arr_VMSME_17_DATA;
  signal VMSME_17_mem_AAAV_dout_nent : t_arr_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSTE_22_mem_A_enb          : t_arr_VMSTE_22_1b;
  signal VMSTE_22_mem_AV_readaddr    : t_arr_VMSTE_22_ADDR;
  signal VMSTE_22_mem_AV_dout        : t_arr_VMSTE_22_DATA;
  signal VMSTE_22_mem_AAV_dout_nent  : t_arr_VMSTE_22_NENT; -- (#page)
  signal VMSTE_16_mem_A_enb          : t_arr_VMSTE_16_1b;
  signal VMSTE_16_mem_AV_readaddr    : t_arr_VMSTE_16_ADDR;
  signal VMSTE_16_mem_AV_dout        : t_arr_VMSTE_16_DATA;
  signal VMSTE_16_mem_AAAV_dout_nent : t_arr_VMSTE_16_NENT; -- (#page)(#bin)
  signal SP_14_mem_A_enb          : t_arr_SP_14_1b;
  signal SP_14_mem_AV_readaddr    : t_arr_SP_14_ADDR;
  signal SP_14_mem_AV_dout        : t_arr_SP_14_DATA;
  signal SP_14_mem_AAV_dout_nent  : t_arr_SP_14_NENT; -- (#page)
  signal TPROJ_60_mem_A_enb          : t_arr_TPROJ_60_1b;
  signal TPROJ_60_mem_AV_readaddr    : t_arr_TPROJ_60_ADDR;
  signal TPROJ_60_mem_AV_dout        : t_arr_TPROJ_60_DATA;
  signal TPROJ_60_mem_AAV_dout_nent  : t_arr_TPROJ_60_NENT; -- (#page)
  signal TPROJ_58_mem_A_enb          : t_arr_TPROJ_58_1b;
  signal TPROJ_58_mem_AV_readaddr    : t_arr_TPROJ_58_ADDR;
  signal TPROJ_58_mem_AV_dout        : t_arr_TPROJ_58_DATA;
  signal TPROJ_58_mem_AAV_dout_nent  : t_arr_TPROJ_58_NENT; -- (#page)
  signal TPAR_70_mem_A_enb          : t_arr_TPAR_70_1b;
  signal TPAR_70_mem_AV_readaddr    : t_arr_TPAR_70_ADDR;
  signal TPAR_70_mem_AV_dout        : t_arr_TPAR_70_DATA;
  signal VMPROJ_24_mem_A_enb          : t_arr_VMPROJ_24_1b;
  signal VMPROJ_24_mem_AV_readaddr    : t_arr_VMPROJ_24_ADDR;
  signal VMPROJ_24_mem_AV_dout        : t_arr_VMPROJ_24_DATA;
  signal VMPROJ_24_mem_AAV_dout_nent  : t_arr_VMPROJ_24_NENT; -- (#page)
  signal AP_60_mem_A_enb          : t_arr_AP_60_1b;
  signal AP_60_mem_AV_readaddr    : t_arr_AP_60_ADDR;
  signal AP_60_mem_AV_dout        : t_arr_AP_60_DATA;
  signal AP_58_mem_A_enb          : t_arr_AP_58_1b;
  signal AP_58_mem_AV_readaddr    : t_arr_AP_58_ADDR;
  signal AP_58_mem_AV_dout        : t_arr_AP_58_DATA;
  signal CM_14_mem_A_enb          : t_arr_CM_14_1b;
  signal CM_14_mem_AV_readaddr    : t_arr_CM_14_ADDR;
  signal CM_14_mem_AV_dout        : t_arr_CM_14_DATA;
  signal CM_14_mem_AAV_dout_nent  : t_arr_CM_14_NENT; -- (#page)
  signal FM_52_mem_A_enb          : t_arr_FM_52_1b;
  signal FM_52_mem_AV_readaddr    : t_arr_FM_52_ADDR;
  signal FM_52_mem_AV_dout        : t_arr_FM_52_DATA;
  signal FM_52_mem_AAV_dout_nent  : t_arr_FM_52_NENT; -- (#page)
  signal VMR_start : std_logic := '0';
  signal TE_start : std_logic := '0';
  signal TC_start : std_logic := '0';
  signal TE_L1PHID14_L2PHIB15_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB15_bendinnertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB15_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB15_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB15_bendoutertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB15_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB16_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB16_bendinnertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB16_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB16_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB16_bendoutertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB16_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB13_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB13_bendinnertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB13_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB13_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB13_bendoutertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB13_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB14_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB14_bendinnertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB14_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB14_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB14_bendoutertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB14_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB15_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB15_bendinnertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB15_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB15_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB15_bendoutertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB15_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB16_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB16_bendinnertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB16_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID15_L2PHIB16_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID15_L2PHIB16_bendoutertable_ce       : std_logic;
  signal TE_L1PHID15_L2PHIB16_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID16_L2PHIB14_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID16_L2PHIB14_bendinnertable_ce       : std_logic;
  signal TE_L1PHID16_L2PHIB14_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID16_L2PHIB14_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID16_L2PHIB14_bendoutertable_ce       : std_logic;
  signal TE_L1PHID16_L2PHIB14_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID16_L2PHIB15_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID16_L2PHIB15_bendinnertable_ce       : std_logic;
  signal TE_L1PHID16_L2PHIB15_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID16_L2PHIB15_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID16_L2PHIB15_bendoutertable_ce       : std_logic;
  signal TE_L1PHID16_L2PHIB15_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID16_L2PHIB16_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID16_L2PHIB16_bendinnertable_ce       : std_logic;
  signal TE_L1PHID16_L2PHIB16_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID16_L2PHIB16_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID16_L2PHIB16_bendoutertable_ce       : std_logic;
  signal TE_L1PHID16_L2PHIB16_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal PR_start : std_logic := '0';
  signal ME_start : std_logic := '0';
  signal MC_start : std_logic := '0';
  signal FT_start : std_logic := '0';

begin

  IL_36_loop : for var in enum_IL_36 generate
  begin

    IL_36 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => IL_36_mem_A_wea(var),
        addra     => IL_36_mem_AV_writeaddr(var),
        dina      => IL_36_mem_AV_din(var),
        clkb      => clk,
        enb       => IL_36_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => IL_36_mem_AV_readaddr(var),
        doutb     => IL_36_mem_AV_dout(var),
        sync_nent => VMR_start,
        nent_o    => IL_36_mem_AAV_dout_nent(var)
      );

  end generate IL_36_loop;


  AS_36_loop : for var in enum_AS_36 generate
  begin

    AS_36 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => AS_36_mem_A_wea(var),
        addra     => AS_36_mem_AV_writeaddr(var),
        dina      => AS_36_mem_AV_din(var),
        clkb      => clk,
        enb       => AS_36_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => AS_36_mem_AV_readaddr(var),
        doutb     => AS_36_mem_AV_dout(var),
        sync_nent => TC_start,
        nent_o    => open
      );

  end generate AS_36_loop;


  VMSME_16_loop : for var in enum_VMSME_16 generate
  begin

    VMSME_16 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => VMSME_16_mem_A_wea(var),
        addra     => VMSME_16_mem_AV_writeaddr(var),
        dina      => VMSME_16_mem_AV_din(var),
        clkb      => clk,
        enb       => VMSME_16_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => VMSME_16_mem_AV_readaddr(var),
        doutb     => VMSME_16_mem_AV_dout(var),
        sync_nent => ME_start,
        nent_o    => VMSME_16_mem_AAAV_dout_nent(var)
      );

  end generate VMSME_16_loop;


  VMSME_17_loop : for var in enum_VMSME_17 generate
  begin

    VMSME_17 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => VMSME_17_mem_A_wea(var),
        addra     => VMSME_17_mem_AV_writeaddr(var),
        dina      => VMSME_17_mem_AV_din(var),
        clkb      => clk,
        enb       => VMSME_17_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => VMSME_17_mem_AV_readaddr(var),
        doutb     => VMSME_17_mem_AV_dout(var),
        sync_nent => ME_start,
        nent_o    => VMSME_17_mem_AAAV_dout_nent(var)
      );

  end generate VMSME_17_loop;


  VMSTE_22_loop : for var in enum_VMSTE_22 generate
  begin

    VMSTE_22 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 22,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => VMSTE_22_mem_A_wea(var),
        addra     => VMSTE_22_mem_AV_writeaddr(var),
        dina      => VMSTE_22_mem_AV_din(var),
        clkb      => clk,
        enb       => VMSTE_22_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => VMSTE_22_mem_AV_readaddr(var),
        doutb     => VMSTE_22_mem_AV_dout(var),
        sync_nent => TE_start,
        nent_o    => VMSTE_22_mem_AAV_dout_nent(var)
      );

  end generate VMSTE_22_loop;


  VMSTE_16_loop : for var in enum_VMSTE_16 generate
  begin

    VMSTE_16 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => VMSTE_16_mem_A_wea(var),
        addra     => VMSTE_16_mem_AV_writeaddr(var),
        dina      => VMSTE_16_mem_AV_din(var),
        clkb      => clk,
        enb       => VMSTE_16_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => VMSTE_16_mem_AV_readaddr(var),
        doutb     => VMSTE_16_mem_AV_dout(var),
        sync_nent => TE_start,
        nent_o    => VMSTE_16_mem_AAAV_dout_nent(var)
      );

  end generate VMSTE_16_loop;


  SP_14_loop : for var in enum_SP_14 generate
  begin

    SP_14 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 14,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => SP_14_mem_A_wea(var),
        addra     => SP_14_mem_AV_writeaddr(var),
        dina      => SP_14_mem_AV_din(var),
        clkb      => clk,
        enb       => SP_14_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => SP_14_mem_AV_readaddr(var),
        doutb     => SP_14_mem_AV_dout(var),
        sync_nent => TC_start,
        nent_o    => SP_14_mem_AAV_dout_nent(var)
      );

  end generate SP_14_loop;


  TPROJ_60_loop : for var in enum_TPROJ_60 generate
  begin

    TPROJ_60 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => TPROJ_60_mem_A_wea(var),
        addra     => TPROJ_60_mem_AV_writeaddr(var),
        dina      => TPROJ_60_mem_AV_din(var),
        clkb      => clk,
        enb       => TPROJ_60_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => TPROJ_60_mem_AV_readaddr(var),
        doutb     => TPROJ_60_mem_AV_dout(var),
        sync_nent => PR_start,
        nent_o    => TPROJ_60_mem_AAV_dout_nent(var)
      );

  end generate TPROJ_60_loop;


  TPROJ_58_loop : for var in enum_TPROJ_58 generate
  begin

    TPROJ_58 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => TPROJ_58_mem_A_wea(var),
        addra     => TPROJ_58_mem_AV_writeaddr(var),
        dina      => TPROJ_58_mem_AV_din(var),
        clkb      => clk,
        enb       => TPROJ_58_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => TPROJ_58_mem_AV_readaddr(var),
        doutb     => TPROJ_58_mem_AV_dout(var),
        sync_nent => PR_start,
        nent_o    => TPROJ_58_mem_AAV_dout_nent(var)
      );

  end generate TPROJ_58_loop;


  TPAR_70_loop : for var in enum_TPAR_70 generate
  begin

    TPAR_70 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 70,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => TPAR_70_mem_A_wea(var),
        addra     => TPAR_70_mem_AV_writeaddr(var),
        dina      => TPAR_70_mem_AV_din(var),
        clkb      => clk,
        enb       => TPAR_70_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => TPAR_70_mem_AV_readaddr(var),
        doutb     => TPAR_70_mem_AV_dout(var),
        sync_nent => FT_start,
        nent_o    => open
      );

  end generate TPAR_70_loop;


  VMPROJ_24_loop : for var in enum_VMPROJ_24 generate
  begin

    VMPROJ_24 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 24,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => VMPROJ_24_mem_A_wea(var),
        addra     => VMPROJ_24_mem_AV_writeaddr(var),
        dina      => VMPROJ_24_mem_AV_din(var),
        clkb      => clk,
        enb       => VMPROJ_24_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => VMPROJ_24_mem_AV_readaddr(var),
        doutb     => VMPROJ_24_mem_AV_dout(var),
        sync_nent => ME_start,
        nent_o    => VMPROJ_24_mem_AAV_dout_nent(var)
      );

  end generate VMPROJ_24_loop;


  AP_60_loop : for var in enum_AP_60 generate
  begin

    AP_60 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => AP_60_mem_A_wea(var),
        addra     => AP_60_mem_AV_writeaddr(var),
        dina      => AP_60_mem_AV_din(var),
        clkb      => clk,
        enb       => AP_60_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => AP_60_mem_AV_readaddr(var),
        doutb     => AP_60_mem_AV_dout(var),
        sync_nent => MC_start,
        nent_o    => open
      );

  end generate AP_60_loop;


  AP_58_loop : for var in enum_AP_58 generate
  begin

    AP_58 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => AP_58_mem_A_wea(var),
        addra     => AP_58_mem_AV_writeaddr(var),
        dina      => AP_58_mem_AV_din(var),
        clkb      => clk,
        enb       => AP_58_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => AP_58_mem_AV_readaddr(var),
        doutb     => AP_58_mem_AV_dout(var),
        sync_nent => MC_start,
        nent_o    => open
      );

  end generate AP_58_loop;


  CM_14_loop : for var in enum_CM_14 generate
  begin

    CM_14 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 14,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => CM_14_mem_A_wea(var),
        addra     => CM_14_mem_AV_writeaddr(var),
        dina      => CM_14_mem_AV_din(var),
        clkb      => clk,
        enb       => CM_14_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => CM_14_mem_AV_readaddr(var),
        doutb     => CM_14_mem_AV_dout(var),
        sync_nent => MC_start,
        nent_o    => CM_14_mem_AAV_dout_nent(var)
      );

  end generate CM_14_loop;


  FM_52_loop : for var in enum_FM_52 generate
  begin

    FM_52 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => FM_52_mem_A_wea(var),
        addra     => FM_52_mem_AV_writeaddr(var),
        dina      => FM_52_mem_AV_din(var),
        clkb      => clk,
        enb       => FM_52_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => FM_52_mem_AV_readaddr(var),
        doutb     => FM_52_mem_AV_dout(var),
        sync_nent => FT_start,
        nent_o    => FM_52_mem_AAV_dout_nent(var)
      );

  end generate FM_52_loop;


  VMR_start <= '1' when IR_done = '1';

  IR_PS10G_1_A : entity work.IR_PS10G_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => IR_done,
      bx_V          => IR_bx_in,
      bx_o_V        => IR_bx_out,
      bx_o_V_ap_vld => IR_bx_out_vld,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS10G_1_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS10G_1_A),
      hInputStubs_V_read     => DL_39_link_read(PS10G_1_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L1PHID_PS10G_1_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L1PHID_PS10G_1_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L1PHID_PS10G_1_A),
      hLinkWord_V => "00100000000000000011",
      hPhBnWord_V => "000000000000"
  );

  IR_PS10G_2_A : entity work.IR_PS10G_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS10G_2_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS10G_2_A),
      hInputStubs_V_read     => DL_39_link_read(PS10G_2_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L1PHID_PS10G_2_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L1PHID_PS10G_2_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L1PHID_PS10G_2_A),
      hLinkWord_V => "00100000000000000011",
      hPhBnWord_V => "000000000000"
  );

  IR_PS10G_2_B : entity work.IR_PS10G_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS10G_2_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS10G_2_B),
      hInputStubs_V_read     => DL_39_link_read(PS10G_2_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L1PHID_PS10G_2_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L1PHID_PS10G_2_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L1PHID_PS10G_2_B),
      hLinkWord_V => "00100000000000000011",
      hPhBnWord_V => "000000000000"
  );

  IR_PS10G_3_A : entity work.IR_PS10G_3_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS10G_3_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS10G_3_A),
      hInputStubs_V_read     => DL_39_link_read(PS10G_3_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L2PHIB_PS10G_3_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L2PHIB_PS10G_3_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L2PHIB_PS10G_3_A),
      hLinkWord_V => "00100000000000000101",
      hPhBnWord_V => "000000000000"
  );

  IR_PS10G_3_B : entity work.IR_PS10G_3_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS10G_3_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS10G_3_B),
      hInputStubs_V_read     => DL_39_link_read(PS10G_3_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L2PHIB_PS10G_3_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L2PHIB_PS10G_3_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L2PHIB_PS10G_3_B),
      hLinkWord_V => "00100000000000000101",
      hPhBnWord_V => "000000000000"
  );

  IR_PS_1_A : entity work.IR_PS_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS_1_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS_1_A),
      hInputStubs_V_read     => DL_39_link_read(PS_1_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L3PHIB_PS_1_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L3PHIB_PS_1_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L3PHIB_PS_1_A),
      hLinkWord_V => "00100000000000000111",
      hPhBnWord_V => "000000000000"
  );

  IR_PS_1_B : entity work.IR_PS_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS_1_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS_1_B),
      hInputStubs_V_read     => DL_39_link_read(PS_1_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L3PHIB_PS_1_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L3PHIB_PS_1_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L3PHIB_PS_1_B),
      hLinkWord_V => "00100000000000000111",
      hPhBnWord_V => "000000000000"
  );

  IR_PS_2_A : entity work.IR_PS_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS_2_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS_2_A),
      hInputStubs_V_read     => DL_39_link_read(PS_2_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L3PHIB_PS_2_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L3PHIB_PS_2_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L3PHIB_PS_2_A),
      hLinkWord_V => "00100000000000000111",
      hPhBnWord_V => "000000000000"
  );

  IR_PS_2_B : entity work.IR_PS_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(PS_2_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(PS_2_B),
      hInputStubs_V_read     => DL_39_link_read(PS_2_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L3PHIB_PS_2_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L3PHIB_PS_2_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L3PHIB_PS_2_B),
      hLinkWord_V => "00100000000000000111",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_1_A : entity work.IR_2S_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_1_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_1_A),
      hInputStubs_V_read     => DL_39_link_read(SS_1_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L4PHIB_2S_1_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L4PHIB_2S_1_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L4PHIB_2S_1_A),
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_36_mem_A_wea(L5PHIB_2S_1_A),
      hOutputStubs_1_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L5PHIB_2S_1_A),
      hOutputStubs_1_dataarray_data_V_d0        => IL_36_mem_AV_din(L5PHIB_2S_1_A),
      hLinkWord_V => "01010000000010111001",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_1_B : entity work.IR_2S_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_1_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_1_B),
      hInputStubs_V_read     => DL_39_link_read(SS_1_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L4PHIB_2S_1_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L4PHIB_2S_1_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L4PHIB_2S_1_B),
      hLinkWord_V => "00110000000000001001",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_2_A : entity work.IR_2S_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_2_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_2_A),
      hInputStubs_V_read     => DL_39_link_read(SS_2_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L5PHIB_2S_2_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L5PHIB_2S_2_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L5PHIB_2S_2_A),
      hLinkWord_V => "00110000000000001011",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_2_B : entity work.IR_2S_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_2_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_2_B),
      hInputStubs_V_read     => DL_39_link_read(SS_2_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L5PHIB_2S_2_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L5PHIB_2S_2_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L5PHIB_2S_2_B),
      hLinkWord_V => "00110000000000001011",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_3_A : entity work.IR_2S_3_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_3_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_3_A),
      hInputStubs_V_read     => DL_39_link_read(SS_3_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L6PHIB_2S_3_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L6PHIB_2S_3_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L6PHIB_2S_3_A),
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_3_B : entity work.IR_2S_3_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_3_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_3_B),
      hInputStubs_V_read     => DL_39_link_read(SS_3_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L6PHIB_2S_3_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L6PHIB_2S_3_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L6PHIB_2S_3_B),
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_4_A : entity work.IR_2S_4_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_4_A),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_4_A),
      hInputStubs_V_read     => DL_39_link_read(SS_4_A),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L6PHIB_2S_4_A),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L6PHIB_2S_4_A),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L6PHIB_2S_4_A),
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "000000000000"
  );

  IR_2S_4_B : entity work.IR_2S_4_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_in,
      hInputStubs_V_dout     => DL_39_link_AV_dout(SS_4_B),
      hInputStubs_V_empty_n  => DL_39_link_empty_neg(SS_4_B),
      hInputStubs_V_read     => DL_39_link_read(SS_4_B),
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_36_mem_A_wea(L6PHIB_2S_4_B),
      hOutputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_writeaddr(L6PHIB_2S_4_B),
      hOutputStubs_0_dataarray_data_V_d0        => IL_36_mem_AV_din(L6PHIB_2S_4_B),
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "000000000000"
  );

  TE_start <= '1' when VMR_done = '1';

  VMR_L1PHID : entity work.VMR_L1PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => VMR_done,
      bx_V          => IR_bx_out,
      bx_o_V        => VMR_bx_out,
      bx_o_V_ap_vld => VMR_bx_out_vld,
      inputStubs_0_dataarray_data_V_ce0       => IL_36_mem_A_enb(L1PHID_PS10G_1_A),
      inputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L1PHID_PS10G_1_A),
      inputStubs_0_dataarray_data_V_q0        => IL_36_mem_AV_dout(L1PHID_PS10G_1_A),
      inputStubs_0_nentries_0_V               => IL_36_mem_AAV_dout_nent(L1PHID_PS10G_1_A)(0),
      inputStubs_0_nentries_1_V               => IL_36_mem_AAV_dout_nent(L1PHID_PS10G_1_A)(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_36_mem_A_enb(L1PHID_PS10G_2_A),
      inputStubs_1_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L1PHID_PS10G_2_A),
      inputStubs_1_dataarray_data_V_q0        => IL_36_mem_AV_dout(L1PHID_PS10G_2_A),
      inputStubs_1_nentries_0_V               => IL_36_mem_AAV_dout_nent(L1PHID_PS10G_2_A)(0),
      inputStubs_1_nentries_1_V               => IL_36_mem_AAV_dout_nent(L1PHID_PS10G_2_A)(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_36_mem_A_enb(L1PHID_PS10G_2_B),
      inputStubs_2_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L1PHID_PS10G_2_B),
      inputStubs_2_dataarray_data_V_q0        => IL_36_mem_AV_dout(L1PHID_PS10G_2_B),
      inputStubs_2_nentries_0_V               => IL_36_mem_AAV_dout_nent(L1PHID_PS10G_2_B)(0),
      inputStubs_2_nentries_1_V               => IL_36_mem_AAV_dout_nent(L1PHID_PS10G_2_B)(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_36_mem_A_wea(L1PHIDn3),
      memoriesAS_0_dataarray_data_V_address0  => AS_36_mem_AV_writeaddr(L1PHIDn3),
      memoriesAS_0_dataarray_data_V_d0        => AS_36_mem_AV_din(L1PHIDn3),
      memoriesTEI_0_0_dataarray_data_V_ce0       => open,
      memoriesTEI_0_0_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID14n4),
      memoriesTEI_0_0_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID14n4),
      memoriesTEI_0_0_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID14n4),
      memoriesTEI_0_1_dataarray_data_V_ce0       => open,
      memoriesTEI_0_1_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID14n5),
      memoriesTEI_0_1_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID14n5),
      memoriesTEI_0_1_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID14n5),
      memoriesTEI_1_0_dataarray_data_V_ce0       => open,
      memoriesTEI_1_0_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID15n1),
      memoriesTEI_1_0_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID15n1),
      memoriesTEI_1_0_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID15n1),
      memoriesTEI_1_1_dataarray_data_V_ce0       => open,
      memoriesTEI_1_1_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID15n2),
      memoriesTEI_1_1_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID15n2),
      memoriesTEI_1_1_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID15n2),
      memoriesTEI_1_2_dataarray_data_V_ce0       => open,
      memoriesTEI_1_2_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID15n3),
      memoriesTEI_1_2_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID15n3),
      memoriesTEI_1_2_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID15n3),
      memoriesTEI_1_3_dataarray_data_V_ce0       => open,
      memoriesTEI_1_3_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID15n4),
      memoriesTEI_1_3_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID15n4),
      memoriesTEI_1_3_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID15n4),
      memoriesTEI_2_0_dataarray_data_V_ce0       => open,
      memoriesTEI_2_0_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID16n1),
      memoriesTEI_2_0_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID16n1),
      memoriesTEI_2_0_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID16n1),
      memoriesTEI_2_1_dataarray_data_V_ce0       => open,
      memoriesTEI_2_1_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID16n2),
      memoriesTEI_2_1_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID16n2),
      memoriesTEI_2_1_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID16n2),
      memoriesTEI_2_2_dataarray_data_V_ce0       => open,
      memoriesTEI_2_2_dataarray_data_V_we0       => VMSTE_22_mem_A_wea(L1PHID16n3),
      memoriesTEI_2_2_dataarray_data_V_address0  => VMSTE_22_mem_AV_writeaddr(L1PHID16n3),
      memoriesTEI_2_2_dataarray_data_V_d0        => VMSTE_22_mem_AV_din(L1PHID16n3)
  );

  VMR_L2PHIB : entity work.VMR_L2PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_out,
      inputStubs_0_dataarray_data_V_ce0       => IL_36_mem_A_enb(L2PHIB_PS10G_3_A),
      inputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L2PHIB_PS10G_3_A),
      inputStubs_0_dataarray_data_V_q0        => IL_36_mem_AV_dout(L2PHIB_PS10G_3_A),
      inputStubs_0_nentries_0_V               => IL_36_mem_AAV_dout_nent(L2PHIB_PS10G_3_A)(0),
      inputStubs_0_nentries_1_V               => IL_36_mem_AAV_dout_nent(L2PHIB_PS10G_3_A)(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_36_mem_A_enb(L2PHIB_PS10G_3_B),
      inputStubs_1_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L2PHIB_PS10G_3_B),
      inputStubs_1_dataarray_data_V_q0        => IL_36_mem_AV_dout(L2PHIB_PS10G_3_B),
      inputStubs_1_nentries_0_V               => IL_36_mem_AAV_dout_nent(L2PHIB_PS10G_3_B)(0),
      inputStubs_1_nentries_1_V               => IL_36_mem_AAV_dout_nent(L2PHIB_PS10G_3_B)(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_36_mem_A_wea(L2PHIBn5),
      memoriesAS_0_dataarray_data_V_address0  => AS_36_mem_AV_writeaddr(L2PHIBn5),
      memoriesAS_0_dataarray_data_V_d0        => AS_36_mem_AV_din(L2PHIBn5),
      memoriesTEO_0_0_dataarray_data_V_ce0       => open,
      memoriesTEO_0_0_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB13n5),
      memoriesTEO_0_0_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB13n5),
      memoriesTEO_0_0_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB13n5),
      memoriesTEO_1_0_dataarray_data_V_ce0       => open,
      memoriesTEO_1_0_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB14n4),
      memoriesTEO_1_0_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB14n4),
      memoriesTEO_1_0_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB14n4),
      memoriesTEO_1_1_dataarray_data_V_ce0       => open,
      memoriesTEO_1_1_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB14n5),
      memoriesTEO_1_1_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB14n5),
      memoriesTEO_1_1_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB14n5),
      memoriesTEO_2_0_dataarray_data_V_ce0       => open,
      memoriesTEO_2_0_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB15n2),
      memoriesTEO_2_0_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB15n2),
      memoriesTEO_2_0_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB15n2),
      memoriesTEO_2_1_dataarray_data_V_ce0       => open,
      memoriesTEO_2_1_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB15n3),
      memoriesTEO_2_1_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB15n3),
      memoriesTEO_2_1_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB15n3),
      memoriesTEO_2_2_dataarray_data_V_ce0       => open,
      memoriesTEO_2_2_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB15n4),
      memoriesTEO_2_2_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB15n4),
      memoriesTEO_2_2_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB15n4),
      memoriesTEO_3_0_dataarray_data_V_ce0       => open,
      memoriesTEO_3_0_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB16n1),
      memoriesTEO_3_0_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB16n1),
      memoriesTEO_3_0_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB16n1),
      memoriesTEO_3_1_dataarray_data_V_ce0       => open,
      memoriesTEO_3_1_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB16n2),
      memoriesTEO_3_1_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB16n2),
      memoriesTEO_3_1_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB16n2),
      memoriesTEO_3_2_dataarray_data_V_ce0       => open,
      memoriesTEO_3_2_dataarray_data_V_we0       => VMSTE_16_mem_A_wea(L2PHIB16n3),
      memoriesTEO_3_2_dataarray_data_V_address0  => VMSTE_16_mem_AV_writeaddr(L2PHIB16n3),
      memoriesTEO_3_2_dataarray_data_V_d0        => VMSTE_16_mem_AV_din(L2PHIB16n3)
  );

  VMR_L3PHIB : entity work.VMR_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_out,
      inputStubs_0_dataarray_data_V_ce0       => IL_36_mem_A_enb(L3PHIB_PS_1_A),
      inputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L3PHIB_PS_1_A),
      inputStubs_0_dataarray_data_V_q0        => IL_36_mem_AV_dout(L3PHIB_PS_1_A),
      inputStubs_0_nentries_0_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_1_A)(0),
      inputStubs_0_nentries_1_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_1_A)(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_36_mem_A_enb(L3PHIB_PS_1_B),
      inputStubs_1_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L3PHIB_PS_1_B),
      inputStubs_1_dataarray_data_V_q0        => IL_36_mem_AV_dout(L3PHIB_PS_1_B),
      inputStubs_1_nentries_0_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_1_B)(0),
      inputStubs_1_nentries_1_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_1_B)(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_36_mem_A_enb(L3PHIB_PS_2_A),
      inputStubs_2_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L3PHIB_PS_2_A),
      inputStubs_2_dataarray_data_V_q0        => IL_36_mem_AV_dout(L3PHIB_PS_2_A),
      inputStubs_2_nentries_0_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_2_A)(0),
      inputStubs_2_nentries_1_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_2_A)(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_36_mem_A_enb(L3PHIB_PS_2_B),
      inputStubs_3_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L3PHIB_PS_2_B),
      inputStubs_3_dataarray_data_V_q0        => IL_36_mem_AV_dout(L3PHIB_PS_2_B),
      inputStubs_3_nentries_0_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_2_B)(0),
      inputStubs_3_nentries_1_V               => IL_36_mem_AAV_dout_nent(L3PHIB_PS_2_B)(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_36_mem_A_wea(L3PHIBn1),
      memoriesAS_0_dataarray_data_V_address0  => AS_36_mem_AV_writeaddr(L3PHIBn1),
      memoriesAS_0_dataarray_data_V_d0        => AS_36_mem_AV_din(L3PHIBn1),
      memoriesME_0_dataarray_data_V_ce0       => open,
      memoriesME_0_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB9n1),
      memoriesME_0_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB9n1),
      memoriesME_0_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB9n1),
      memoriesME_1_dataarray_data_V_ce0       => open,
      memoriesME_1_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB10n1),
      memoriesME_1_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB10n1),
      memoriesME_1_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB10n1),
      memoriesME_2_dataarray_data_V_ce0       => open,
      memoriesME_2_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB11n1),
      memoriesME_2_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB11n1),
      memoriesME_2_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB11n1),
      memoriesME_3_dataarray_data_V_ce0       => open,
      memoriesME_3_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB12n1),
      memoriesME_3_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB12n1),
      memoriesME_3_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB12n1),
      memoriesME_4_dataarray_data_V_ce0       => open,
      memoriesME_4_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB13n1),
      memoriesME_4_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB13n1),
      memoriesME_4_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB13n1),
      memoriesME_5_dataarray_data_V_ce0       => open,
      memoriesME_5_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB14n1),
      memoriesME_5_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB14n1),
      memoriesME_5_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB14n1),
      memoriesME_6_dataarray_data_V_ce0       => open,
      memoriesME_6_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB15n1),
      memoriesME_6_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB15n1),
      memoriesME_6_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB15n1),
      memoriesME_7_dataarray_data_V_ce0       => open,
      memoriesME_7_dataarray_data_V_we0       => VMSME_16_mem_A_wea(L3PHIB16n1),
      memoriesME_7_dataarray_data_V_address0  => VMSME_16_mem_AV_writeaddr(L3PHIB16n1),
      memoriesME_7_dataarray_data_V_d0        => VMSME_16_mem_AV_din(L3PHIB16n1)
  );

  VMR_L4PHIB : entity work.VMR_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_out,
      inputStubs_0_dataarray_data_V_ce0       => IL_36_mem_A_enb(L4PHIB_2S_1_A),
      inputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L4PHIB_2S_1_A),
      inputStubs_0_dataarray_data_V_q0        => IL_36_mem_AV_dout(L4PHIB_2S_1_A),
      inputStubs_0_nentries_0_V               => IL_36_mem_AAV_dout_nent(L4PHIB_2S_1_A)(0),
      inputStubs_0_nentries_1_V               => IL_36_mem_AAV_dout_nent(L4PHIB_2S_1_A)(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_36_mem_A_enb(L4PHIB_2S_1_B),
      inputStubs_1_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L4PHIB_2S_1_B),
      inputStubs_1_dataarray_data_V_q0        => IL_36_mem_AV_dout(L4PHIB_2S_1_B),
      inputStubs_1_nentries_0_V               => IL_36_mem_AAV_dout_nent(L4PHIB_2S_1_B)(0),
      inputStubs_1_nentries_1_V               => IL_36_mem_AAV_dout_nent(L4PHIB_2S_1_B)(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_36_mem_A_wea(L4PHIBn1),
      memoriesAS_0_dataarray_data_V_address0  => AS_36_mem_AV_writeaddr(L4PHIBn1),
      memoriesAS_0_dataarray_data_V_d0        => AS_36_mem_AV_din(L4PHIBn1),
      memoriesME_0_dataarray_data_V_ce0       => open,
      memoriesME_0_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB9n1),
      memoriesME_0_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB9n1),
      memoriesME_0_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB9n1),
      memoriesME_1_dataarray_data_V_ce0       => open,
      memoriesME_1_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB10n1),
      memoriesME_1_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB10n1),
      memoriesME_1_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB10n1),
      memoriesME_2_dataarray_data_V_ce0       => open,
      memoriesME_2_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB11n1),
      memoriesME_2_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB11n1),
      memoriesME_2_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB11n1),
      memoriesME_3_dataarray_data_V_ce0       => open,
      memoriesME_3_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB12n1),
      memoriesME_3_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB12n1),
      memoriesME_3_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB12n1),
      memoriesME_4_dataarray_data_V_ce0       => open,
      memoriesME_4_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB13n1),
      memoriesME_4_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB13n1),
      memoriesME_4_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB13n1),
      memoriesME_5_dataarray_data_V_ce0       => open,
      memoriesME_5_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB14n1),
      memoriesME_5_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB14n1),
      memoriesME_5_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB14n1),
      memoriesME_6_dataarray_data_V_ce0       => open,
      memoriesME_6_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB15n1),
      memoriesME_6_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB15n1),
      memoriesME_6_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB15n1),
      memoriesME_7_dataarray_data_V_ce0       => open,
      memoriesME_7_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L4PHIB16n1),
      memoriesME_7_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L4PHIB16n1),
      memoriesME_7_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L4PHIB16n1)
  );

  VMR_L5PHIB : entity work.VMR_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_out,
      inputStubs_0_dataarray_data_V_ce0       => IL_36_mem_A_enb(L5PHIB_2S_1_A),
      inputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L5PHIB_2S_1_A),
      inputStubs_0_dataarray_data_V_q0        => IL_36_mem_AV_dout(L5PHIB_2S_1_A),
      inputStubs_0_nentries_0_V               => IL_36_mem_AAV_dout_nent(L5PHIB_2S_1_A)(0),
      inputStubs_0_nentries_1_V               => IL_36_mem_AAV_dout_nent(L5PHIB_2S_1_A)(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_36_mem_A_enb(L5PHIB_2S_2_A),
      inputStubs_1_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L5PHIB_2S_2_A),
      inputStubs_1_dataarray_data_V_q0        => IL_36_mem_AV_dout(L5PHIB_2S_2_A),
      inputStubs_1_nentries_0_V               => IL_36_mem_AAV_dout_nent(L5PHIB_2S_2_A)(0),
      inputStubs_1_nentries_1_V               => IL_36_mem_AAV_dout_nent(L5PHIB_2S_2_A)(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_36_mem_A_enb(L5PHIB_2S_2_B),
      inputStubs_2_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L5PHIB_2S_2_B),
      inputStubs_2_dataarray_data_V_q0        => IL_36_mem_AV_dout(L5PHIB_2S_2_B),
      inputStubs_2_nentries_0_V               => IL_36_mem_AAV_dout_nent(L5PHIB_2S_2_B)(0),
      inputStubs_2_nentries_1_V               => IL_36_mem_AAV_dout_nent(L5PHIB_2S_2_B)(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_36_mem_A_wea(L5PHIBn1),
      memoriesAS_0_dataarray_data_V_address0  => AS_36_mem_AV_writeaddr(L5PHIBn1),
      memoriesAS_0_dataarray_data_V_d0        => AS_36_mem_AV_din(L5PHIBn1),
      memoriesME_0_dataarray_data_V_ce0       => open,
      memoriesME_0_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB9n1),
      memoriesME_0_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB9n1),
      memoriesME_0_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB9n1),
      memoriesME_1_dataarray_data_V_ce0       => open,
      memoriesME_1_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB10n1),
      memoriesME_1_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB10n1),
      memoriesME_1_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB10n1),
      memoriesME_2_dataarray_data_V_ce0       => open,
      memoriesME_2_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB11n1),
      memoriesME_2_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB11n1),
      memoriesME_2_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB11n1),
      memoriesME_3_dataarray_data_V_ce0       => open,
      memoriesME_3_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB12n1),
      memoriesME_3_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB12n1),
      memoriesME_3_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB12n1),
      memoriesME_4_dataarray_data_V_ce0       => open,
      memoriesME_4_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB13n1),
      memoriesME_4_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB13n1),
      memoriesME_4_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB13n1),
      memoriesME_5_dataarray_data_V_ce0       => open,
      memoriesME_5_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB14n1),
      memoriesME_5_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB14n1),
      memoriesME_5_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB14n1),
      memoriesME_6_dataarray_data_V_ce0       => open,
      memoriesME_6_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB15n1),
      memoriesME_6_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB15n1),
      memoriesME_6_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB15n1),
      memoriesME_7_dataarray_data_V_ce0       => open,
      memoriesME_7_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L5PHIB16n1),
      memoriesME_7_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L5PHIB16n1),
      memoriesME_7_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L5PHIB16n1)
  );

  VMR_L6PHIB : entity work.VMR_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_bx_out,
      inputStubs_0_dataarray_data_V_ce0       => IL_36_mem_A_enb(L6PHIB_2S_3_A),
      inputStubs_0_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L6PHIB_2S_3_A),
      inputStubs_0_dataarray_data_V_q0        => IL_36_mem_AV_dout(L6PHIB_2S_3_A),
      inputStubs_0_nentries_0_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_3_A)(0),
      inputStubs_0_nentries_1_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_3_A)(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_36_mem_A_enb(L6PHIB_2S_3_B),
      inputStubs_1_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L6PHIB_2S_3_B),
      inputStubs_1_dataarray_data_V_q0        => IL_36_mem_AV_dout(L6PHIB_2S_3_B),
      inputStubs_1_nentries_0_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_3_B)(0),
      inputStubs_1_nentries_1_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_3_B)(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_36_mem_A_enb(L6PHIB_2S_4_A),
      inputStubs_2_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L6PHIB_2S_4_A),
      inputStubs_2_dataarray_data_V_q0        => IL_36_mem_AV_dout(L6PHIB_2S_4_A),
      inputStubs_2_nentries_0_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_4_A)(0),
      inputStubs_2_nentries_1_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_4_A)(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_36_mem_A_enb(L6PHIB_2S_4_B),
      inputStubs_3_dataarray_data_V_address0  => IL_36_mem_AV_readaddr(L6PHIB_2S_4_B),
      inputStubs_3_dataarray_data_V_q0        => IL_36_mem_AV_dout(L6PHIB_2S_4_B),
      inputStubs_3_nentries_0_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_4_B)(0),
      inputStubs_3_nentries_1_V               => IL_36_mem_AAV_dout_nent(L6PHIB_2S_4_B)(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_36_mem_A_wea(L6PHIBn1),
      memoriesAS_0_dataarray_data_V_address0  => AS_36_mem_AV_writeaddr(L6PHIBn1),
      memoriesAS_0_dataarray_data_V_d0        => AS_36_mem_AV_din(L6PHIBn1),
      memoriesME_0_dataarray_data_V_ce0       => open,
      memoriesME_0_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB9n1),
      memoriesME_0_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB9n1),
      memoriesME_0_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB9n1),
      memoriesME_1_dataarray_data_V_ce0       => open,
      memoriesME_1_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB10n1),
      memoriesME_1_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB10n1),
      memoriesME_1_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB10n1),
      memoriesME_2_dataarray_data_V_ce0       => open,
      memoriesME_2_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB11n1),
      memoriesME_2_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB11n1),
      memoriesME_2_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB11n1),
      memoriesME_3_dataarray_data_V_ce0       => open,
      memoriesME_3_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB12n1),
      memoriesME_3_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB12n1),
      memoriesME_3_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB12n1),
      memoriesME_4_dataarray_data_V_ce0       => open,
      memoriesME_4_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB13n1),
      memoriesME_4_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB13n1),
      memoriesME_4_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB13n1),
      memoriesME_5_dataarray_data_V_ce0       => open,
      memoriesME_5_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB14n1),
      memoriesME_5_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB14n1),
      memoriesME_5_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB14n1),
      memoriesME_6_dataarray_data_V_ce0       => open,
      memoriesME_6_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB15n1),
      memoriesME_6_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB15n1),
      memoriesME_6_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB15n1),
      memoriesME_7_dataarray_data_V_ce0       => open,
      memoriesME_7_dataarray_data_V_we0       => VMSME_17_mem_A_wea(L6PHIB16n1),
      memoriesME_7_dataarray_data_V_address0  => VMSME_17_mem_AV_writeaddr(L6PHIB16n1),
      memoriesME_7_dataarray_data_V_d0        => VMSME_17_mem_AV_din(L6PHIB16n1)
  );


  TE_L1PHID14_L2PHIB15_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID14_L2PHIB15_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB15_bendinnertable_addr,
      ce        => TE_L1PHID14_L2PHIB15_bendinnertable_ce,
      dout      => TE_L1PHID14_L2PHIB15_bendinnertable_dout
  );


  TE_L1PHID14_L2PHIB15_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID14_L2PHIB15_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB15_bendoutertable_addr,
      ce        => TE_L1PHID14_L2PHIB15_bendoutertable_ce,
      dout      => TE_L1PHID14_L2PHIB15_bendoutertable_dout
  );

  TC_start <= '1' when TE_done = '1';

  TE_L1PHID14_L2PHIB15 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => TE_done,
      bx_V          => VMR_bx_out,
      bx_o_V        => TE_bx_out,
      bx_o_V_ap_vld => TE_bx_out_vld,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID14n4),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID14n4),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID14n4),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n4)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n4)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB15n2),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB15n2),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB15n2),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n2)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID14_L2PHIB15_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID14_L2PHIB15_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID14_L2PHIB15_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID14_L2PHIB15_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID14_L2PHIB15_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID14_L2PHIB15_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID14_L2PHIB15),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID14_L2PHIB15),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID14_L2PHIB15)
  );


  TE_L1PHID14_L2PHIB16_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID14_L2PHIB16_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB16_bendinnertable_addr,
      ce        => TE_L1PHID14_L2PHIB16_bendinnertable_ce,
      dout      => TE_L1PHID14_L2PHIB16_bendinnertable_dout
  );


  TE_L1PHID14_L2PHIB16_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID14_L2PHIB16_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB16_bendoutertable_addr,
      ce        => TE_L1PHID14_L2PHIB16_bendoutertable_ce,
      dout      => TE_L1PHID14_L2PHIB16_bendoutertable_dout
  );

  TE_L1PHID14_L2PHIB16 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID14n5),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID14n5),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID14n5),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n5)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n5)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB16n1),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB16n1),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB16n1),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n1)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID14_L2PHIB16_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID14_L2PHIB16_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID14_L2PHIB16_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID14_L2PHIB16_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID14_L2PHIB16_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID14_L2PHIB16_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID14_L2PHIB16),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID14_L2PHIB16),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID14_L2PHIB16)
  );


  TE_L1PHID15_L2PHIB13_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB13_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB13_bendinnertable_addr,
      ce        => TE_L1PHID15_L2PHIB13_bendinnertable_ce,
      dout      => TE_L1PHID15_L2PHIB13_bendinnertable_dout
  );


  TE_L1PHID15_L2PHIB13_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB13_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB13_bendoutertable_addr,
      ce        => TE_L1PHID15_L2PHIB13_bendoutertable_ce,
      dout      => TE_L1PHID15_L2PHIB13_bendoutertable_dout
  );

  TE_L1PHID15_L2PHIB13 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID15n1),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID15n1),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID15n1),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n1)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n1)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB13n5),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB13n5),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB13n5),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n5)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID15_L2PHIB13_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID15_L2PHIB13_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID15_L2PHIB13_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID15_L2PHIB13_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID15_L2PHIB13_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID15_L2PHIB13_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID15_L2PHIB13),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID15_L2PHIB13),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID15_L2PHIB13)
  );


  TE_L1PHID15_L2PHIB14_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB14_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB14_bendinnertable_addr,
      ce        => TE_L1PHID15_L2PHIB14_bendinnertable_ce,
      dout      => TE_L1PHID15_L2PHIB14_bendinnertable_dout
  );


  TE_L1PHID15_L2PHIB14_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB14_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB14_bendoutertable_addr,
      ce        => TE_L1PHID15_L2PHIB14_bendoutertable_ce,
      dout      => TE_L1PHID15_L2PHIB14_bendoutertable_dout
  );

  TE_L1PHID15_L2PHIB14 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID15n2),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID15n2),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID15n2),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n2)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n2)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB14n4),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB14n4),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB14n4),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n4)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID15_L2PHIB14_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID15_L2PHIB14_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID15_L2PHIB14_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID15_L2PHIB14_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID15_L2PHIB14_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID15_L2PHIB14_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID15_L2PHIB14),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID15_L2PHIB14),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID15_L2PHIB14)
  );


  TE_L1PHID15_L2PHIB15_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB15_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB15_bendinnertable_addr,
      ce        => TE_L1PHID15_L2PHIB15_bendinnertable_ce,
      dout      => TE_L1PHID15_L2PHIB15_bendinnertable_dout
  );


  TE_L1PHID15_L2PHIB15_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB15_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB15_bendoutertable_addr,
      ce        => TE_L1PHID15_L2PHIB15_bendoutertable_ce,
      dout      => TE_L1PHID15_L2PHIB15_bendoutertable_dout
  );

  TE_L1PHID15_L2PHIB15 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID15n3),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID15n3),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID15n3),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n3)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n3)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB15n3),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB15n3),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB15n3),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n3)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID15_L2PHIB15_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID15_L2PHIB15_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID15_L2PHIB15_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID15_L2PHIB15_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID15_L2PHIB15_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID15_L2PHIB15_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID15_L2PHIB15),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID15_L2PHIB15),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID15_L2PHIB15)
  );


  TE_L1PHID15_L2PHIB16_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB16_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB16_bendinnertable_addr,
      ce        => TE_L1PHID15_L2PHIB16_bendinnertable_ce,
      dout      => TE_L1PHID15_L2PHIB16_bendinnertable_dout
  );


  TE_L1PHID15_L2PHIB16_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID15_L2PHIB16_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID15_L2PHIB16_bendoutertable_addr,
      ce        => TE_L1PHID15_L2PHIB16_bendoutertable_ce,
      dout      => TE_L1PHID15_L2PHIB16_bendoutertable_dout
  );

  TE_L1PHID15_L2PHIB16 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID15n4),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID15n4),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID15n4),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n4)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID15n4)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB16n2),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB16n2),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB16n2),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n2)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID15_L2PHIB16_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID15_L2PHIB16_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID15_L2PHIB16_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID15_L2PHIB16_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID15_L2PHIB16_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID15_L2PHIB16_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID15_L2PHIB16),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID15_L2PHIB16),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID15_L2PHIB16)
  );


  TE_L1PHID16_L2PHIB14_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID16_L2PHIB14_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID16_L2PHIB14_bendinnertable_addr,
      ce        => TE_L1PHID16_L2PHIB14_bendinnertable_ce,
      dout      => TE_L1PHID16_L2PHIB14_bendinnertable_dout
  );


  TE_L1PHID16_L2PHIB14_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID16_L2PHIB14_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID16_L2PHIB14_bendoutertable_addr,
      ce        => TE_L1PHID16_L2PHIB14_bendoutertable_ce,
      dout      => TE_L1PHID16_L2PHIB14_bendoutertable_dout
  );

  TE_L1PHID16_L2PHIB14 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID16n1),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID16n1),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID16n1),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID16n1)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID16n1)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB14n5),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB14n5),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB14n5),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n5)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID16_L2PHIB14_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID16_L2PHIB14_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID16_L2PHIB14_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID16_L2PHIB14_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID16_L2PHIB14_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID16_L2PHIB14_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID16_L2PHIB14),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID16_L2PHIB14),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID16_L2PHIB14)
  );


  TE_L1PHID16_L2PHIB15_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID16_L2PHIB15_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID16_L2PHIB15_bendinnertable_addr,
      ce        => TE_L1PHID16_L2PHIB15_bendinnertable_ce,
      dout      => TE_L1PHID16_L2PHIB15_bendinnertable_dout
  );


  TE_L1PHID16_L2PHIB15_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID16_L2PHIB15_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID16_L2PHIB15_bendoutertable_addr,
      ce        => TE_L1PHID16_L2PHIB15_bendoutertable_ce,
      dout      => TE_L1PHID16_L2PHIB15_bendoutertable_dout
  );

  TE_L1PHID16_L2PHIB15 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID16n2),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID16n2),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID16n2),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID16n2)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID16n2)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB15n4),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB15n4),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB15n4),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n4)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID16_L2PHIB15_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID16_L2PHIB15_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID16_L2PHIB15_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID16_L2PHIB15_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID16_L2PHIB15_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID16_L2PHIB15_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID16_L2PHIB15),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID16_L2PHIB15),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID16_L2PHIB15)
  );


  TE_L1PHID16_L2PHIB16_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID16_L2PHIB16_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID16_L2PHIB16_bendinnertable_addr,
      ce        => TE_L1PHID16_L2PHIB16_bendinnertable_ce,
      dout      => TE_L1PHID16_L2PHIB16_bendinnertable_dout
  );


  TE_L1PHID16_L2PHIB16_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => getDirEMDATA & "LUTs/TE_L1PHID16_L2PHIB16_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID16_L2PHIB16_bendoutertable_addr,
      ce        => TE_L1PHID16_L2PHIB16_bendoutertable_ce,
      dout      => TE_L1PHID16_L2PHIB16_bendoutertable_dout
  );

  TE_L1PHID16_L2PHIB16 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_bx_out,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID16n3),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID16n3),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID16n3),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID16n3)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID16n3)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB16n3),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB16n3),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB16n3),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB16n3)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID16_L2PHIB16_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID16_L2PHIB16_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID16_L2PHIB16_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID16_L2PHIB16_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID16_L2PHIB16_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID16_L2PHIB16_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID16_L2PHIB16),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID16_L2PHIB16),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID16_L2PHIB16)
  );

  PR_start <= '1' when TC_done = '1';

  TC_L1L2F : entity work.TC_L1L2F
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => TC_done,
      bx_V          => TE_bx_out,
      bx_o_V        => TC_bx_out,
      bx_o_V_ap_vld => TC_bx_out_vld,
      innerStubs_0_dataarray_data_V_ce0       => AS_36_mem_A_enb(L1PHIDn3),
      innerStubs_0_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L1PHIDn3),
      innerStubs_0_dataarray_data_V_q0        => AS_36_mem_AV_dout(L1PHIDn3),
      outerStubs_0_dataarray_data_V_ce0       => AS_36_mem_A_enb(L2PHIBn5),
      outerStubs_0_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L2PHIBn5),
      outerStubs_0_dataarray_data_V_q0        => AS_36_mem_AV_dout(L2PHIBn5),
      stubPairs_0_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID14_L2PHIB15),
      stubPairs_0_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID14_L2PHIB15),
      stubPairs_0_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID14_L2PHIB15),
      stubPairs_0_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB15)(0),
      stubPairs_0_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB15)(1),
      stubPairs_1_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID14_L2PHIB16),
      stubPairs_1_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID14_L2PHIB16),
      stubPairs_1_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID14_L2PHIB16),
      stubPairs_1_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB16)(0),
      stubPairs_1_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB16)(1),
      stubPairs_2_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID15_L2PHIB13),
      stubPairs_2_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID15_L2PHIB13),
      stubPairs_2_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID15_L2PHIB13),
      stubPairs_2_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB13)(0),
      stubPairs_2_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB13)(1),
      stubPairs_3_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID15_L2PHIB14),
      stubPairs_3_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID15_L2PHIB14),
      stubPairs_3_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID15_L2PHIB14),
      stubPairs_3_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB14)(0),
      stubPairs_3_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB14)(1),
      stubPairs_4_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID15_L2PHIB15),
      stubPairs_4_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID15_L2PHIB15),
      stubPairs_4_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID15_L2PHIB15),
      stubPairs_4_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB15)(0),
      stubPairs_4_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB15)(1),
      stubPairs_5_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID15_L2PHIB16),
      stubPairs_5_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID15_L2PHIB16),
      stubPairs_5_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID15_L2PHIB16),
      stubPairs_5_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB16)(0),
      stubPairs_5_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID15_L2PHIB16)(1),
      stubPairs_6_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID16_L2PHIB14),
      stubPairs_6_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID16_L2PHIB14),
      stubPairs_6_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID16_L2PHIB14),
      stubPairs_6_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID16_L2PHIB14)(0),
      stubPairs_6_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID16_L2PHIB14)(1),
      stubPairs_7_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID16_L2PHIB15),
      stubPairs_7_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID16_L2PHIB15),
      stubPairs_7_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID16_L2PHIB15),
      stubPairs_7_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID16_L2PHIB15)(0),
      stubPairs_7_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID16_L2PHIB15)(1),
      stubPairs_8_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID16_L2PHIB16),
      stubPairs_8_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID16_L2PHIB16),
      stubPairs_8_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID16_L2PHIB16),
      stubPairs_8_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID16_L2PHIB16)(0),
      stubPairs_8_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID16_L2PHIB16)(1),
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_70_mem_A_wea(L1L2F),
      trackletParameters_dataarray_data_V_address0  => TPAR_70_mem_AV_writeaddr(L1L2F),
      trackletParameters_dataarray_data_V_d0        => TPAR_70_mem_AV_din(L1L2F),
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => TPROJ_60_mem_A_wea(L1L2F_L3PHIB),
      projout_barrel_ps_13_dataarray_data_V_address0  => TPROJ_60_mem_AV_writeaddr(L1L2F_L3PHIB),
      projout_barrel_ps_13_dataarray_data_V_d0        => TPROJ_60_mem_AV_din(L1L2F_L3PHIB),
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2F_L4PHIB),
      projout_barrel_2s_1_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2F_L4PHIB),
      projout_barrel_2s_1_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2F_L4PHIB),
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2F_L5PHIB),
      projout_barrel_2s_5_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2F_L5PHIB),
      projout_barrel_2s_5_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2F_L5PHIB),
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2F_L6PHIB),
      projout_barrel_2s_9_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2F_L6PHIB),
      projout_barrel_2s_9_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2F_L6PHIB)
  );

  ME_start <= '1' when PR_done = '1';

  PR_L3PHIB : entity work.PR_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => PR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => PR_done,
      bx_V          => TC_bx_out,
      bx_o_V        => PR_bx_out,
      bx_o_V_ap_vld => PR_bx_out_vld,
      projin_0_dataarray_data_V_ce0       => TPROJ_60_mem_A_enb(L1L2F_L3PHIB),
      projin_0_dataarray_data_V_address0  => TPROJ_60_mem_AV_readaddr(L1L2F_L3PHIB),
      projin_0_dataarray_data_V_q0        => TPROJ_60_mem_AV_dout(L1L2F_L3PHIB),
      projin_0_nentries_0_V               => TPROJ_60_mem_AAV_dout_nent(L1L2F_L3PHIB)(0),
      projin_0_nentries_1_V               => TPROJ_60_mem_AAV_dout_nent(L1L2F_L3PHIB)(1),
      allprojout_dataarray_data_V_ce0       => open,
      allprojout_dataarray_data_V_we0       => AP_60_mem_A_wea(L3PHIB),
      allprojout_dataarray_data_V_address0  => AP_60_mem_AV_writeaddr(L3PHIB),
      allprojout_dataarray_data_V_d0        => AP_60_mem_AV_din(L3PHIB),
      vmprojout_0_dataarray_data_V_ce0       => open,
      vmprojout_0_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB9),
      vmprojout_0_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB9),
      vmprojout_0_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB9),
      vmprojout_1_dataarray_data_V_ce0       => open,
      vmprojout_1_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB10),
      vmprojout_1_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB10),
      vmprojout_1_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB10),
      vmprojout_2_dataarray_data_V_ce0       => open,
      vmprojout_2_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB11),
      vmprojout_2_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB11),
      vmprojout_2_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB11),
      vmprojout_3_dataarray_data_V_ce0       => open,
      vmprojout_3_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB12),
      vmprojout_3_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB12),
      vmprojout_3_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB12),
      vmprojout_4_dataarray_data_V_ce0       => open,
      vmprojout_4_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB13),
      vmprojout_4_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB13),
      vmprojout_4_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB13),
      vmprojout_5_dataarray_data_V_ce0       => open,
      vmprojout_5_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB14),
      vmprojout_5_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB14),
      vmprojout_5_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB14),
      vmprojout_6_dataarray_data_V_ce0       => open,
      vmprojout_6_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB15),
      vmprojout_6_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB15),
      vmprojout_6_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB15),
      vmprojout_7_dataarray_data_V_ce0       => open,
      vmprojout_7_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L3PHIB16),
      vmprojout_7_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L3PHIB16),
      vmprojout_7_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L3PHIB16)
  );

  PR_L4PHIB : entity work.PR_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => PR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TC_bx_out,
      projin_0_dataarray_data_V_ce0       => TPROJ_58_mem_A_enb(L1L2F_L4PHIB),
      projin_0_dataarray_data_V_address0  => TPROJ_58_mem_AV_readaddr(L1L2F_L4PHIB),
      projin_0_dataarray_data_V_q0        => TPROJ_58_mem_AV_dout(L1L2F_L4PHIB),
      projin_0_nentries_0_V               => TPROJ_58_mem_AAV_dout_nent(L1L2F_L4PHIB)(0),
      projin_0_nentries_1_V               => TPROJ_58_mem_AAV_dout_nent(L1L2F_L4PHIB)(1),
      allprojout_dataarray_data_V_ce0       => open,
      allprojout_dataarray_data_V_we0       => AP_58_mem_A_wea(L4PHIB),
      allprojout_dataarray_data_V_address0  => AP_58_mem_AV_writeaddr(L4PHIB),
      allprojout_dataarray_data_V_d0        => AP_58_mem_AV_din(L4PHIB),
      vmprojout_0_dataarray_data_V_ce0       => open,
      vmprojout_0_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB9),
      vmprojout_0_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB9),
      vmprojout_0_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB9),
      vmprojout_1_dataarray_data_V_ce0       => open,
      vmprojout_1_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB10),
      vmprojout_1_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB10),
      vmprojout_1_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB10),
      vmprojout_2_dataarray_data_V_ce0       => open,
      vmprojout_2_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB11),
      vmprojout_2_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB11),
      vmprojout_2_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB11),
      vmprojout_3_dataarray_data_V_ce0       => open,
      vmprojout_3_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB12),
      vmprojout_3_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB12),
      vmprojout_3_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB12),
      vmprojout_4_dataarray_data_V_ce0       => open,
      vmprojout_4_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB13),
      vmprojout_4_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB13),
      vmprojout_4_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB13),
      vmprojout_5_dataarray_data_V_ce0       => open,
      vmprojout_5_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB14),
      vmprojout_5_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB14),
      vmprojout_5_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB14),
      vmprojout_6_dataarray_data_V_ce0       => open,
      vmprojout_6_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB15),
      vmprojout_6_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB15),
      vmprojout_6_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB15),
      vmprojout_7_dataarray_data_V_ce0       => open,
      vmprojout_7_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L4PHIB16),
      vmprojout_7_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L4PHIB16),
      vmprojout_7_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L4PHIB16)
  );

  PR_L5PHIB : entity work.PR_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => PR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TC_bx_out,
      projin_0_dataarray_data_V_ce0       => TPROJ_58_mem_A_enb(L1L2F_L5PHIB),
      projin_0_dataarray_data_V_address0  => TPROJ_58_mem_AV_readaddr(L1L2F_L5PHIB),
      projin_0_dataarray_data_V_q0        => TPROJ_58_mem_AV_dout(L1L2F_L5PHIB),
      projin_0_nentries_0_V               => TPROJ_58_mem_AAV_dout_nent(L1L2F_L5PHIB)(0),
      projin_0_nentries_1_V               => TPROJ_58_mem_AAV_dout_nent(L1L2F_L5PHIB)(1),
      allprojout_dataarray_data_V_ce0       => open,
      allprojout_dataarray_data_V_we0       => AP_58_mem_A_wea(L5PHIB),
      allprojout_dataarray_data_V_address0  => AP_58_mem_AV_writeaddr(L5PHIB),
      allprojout_dataarray_data_V_d0        => AP_58_mem_AV_din(L5PHIB),
      vmprojout_0_dataarray_data_V_ce0       => open,
      vmprojout_0_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB9),
      vmprojout_0_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB9),
      vmprojout_0_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB9),
      vmprojout_1_dataarray_data_V_ce0       => open,
      vmprojout_1_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB10),
      vmprojout_1_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB10),
      vmprojout_1_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB10),
      vmprojout_2_dataarray_data_V_ce0       => open,
      vmprojout_2_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB11),
      vmprojout_2_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB11),
      vmprojout_2_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB11),
      vmprojout_3_dataarray_data_V_ce0       => open,
      vmprojout_3_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB12),
      vmprojout_3_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB12),
      vmprojout_3_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB12),
      vmprojout_4_dataarray_data_V_ce0       => open,
      vmprojout_4_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB13),
      vmprojout_4_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB13),
      vmprojout_4_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB13),
      vmprojout_5_dataarray_data_V_ce0       => open,
      vmprojout_5_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB14),
      vmprojout_5_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB14),
      vmprojout_5_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB14),
      vmprojout_6_dataarray_data_V_ce0       => open,
      vmprojout_6_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB15),
      vmprojout_6_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB15),
      vmprojout_6_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB15),
      vmprojout_7_dataarray_data_V_ce0       => open,
      vmprojout_7_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L5PHIB16),
      vmprojout_7_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L5PHIB16),
      vmprojout_7_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L5PHIB16)
  );

  PR_L6PHIB : entity work.PR_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => PR_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TC_bx_out,
      projin_0_dataarray_data_V_ce0       => TPROJ_58_mem_A_enb(L1L2F_L6PHIB),
      projin_0_dataarray_data_V_address0  => TPROJ_58_mem_AV_readaddr(L1L2F_L6PHIB),
      projin_0_dataarray_data_V_q0        => TPROJ_58_mem_AV_dout(L1L2F_L6PHIB),
      projin_0_nentries_0_V               => TPROJ_58_mem_AAV_dout_nent(L1L2F_L6PHIB)(0),
      projin_0_nentries_1_V               => TPROJ_58_mem_AAV_dout_nent(L1L2F_L6PHIB)(1),
      allprojout_dataarray_data_V_ce0       => open,
      allprojout_dataarray_data_V_we0       => AP_58_mem_A_wea(L6PHIB),
      allprojout_dataarray_data_V_address0  => AP_58_mem_AV_writeaddr(L6PHIB),
      allprojout_dataarray_data_V_d0        => AP_58_mem_AV_din(L6PHIB),
      vmprojout_0_dataarray_data_V_ce0       => open,
      vmprojout_0_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB9),
      vmprojout_0_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB9),
      vmprojout_0_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB9),
      vmprojout_1_dataarray_data_V_ce0       => open,
      vmprojout_1_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB10),
      vmprojout_1_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB10),
      vmprojout_1_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB10),
      vmprojout_2_dataarray_data_V_ce0       => open,
      vmprojout_2_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB11),
      vmprojout_2_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB11),
      vmprojout_2_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB11),
      vmprojout_3_dataarray_data_V_ce0       => open,
      vmprojout_3_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB12),
      vmprojout_3_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB12),
      vmprojout_3_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB12),
      vmprojout_4_dataarray_data_V_ce0       => open,
      vmprojout_4_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB13),
      vmprojout_4_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB13),
      vmprojout_4_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB13),
      vmprojout_5_dataarray_data_V_ce0       => open,
      vmprojout_5_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB14),
      vmprojout_5_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB14),
      vmprojout_5_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB14),
      vmprojout_6_dataarray_data_V_ce0       => open,
      vmprojout_6_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB15),
      vmprojout_6_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB15),
      vmprojout_6_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB15),
      vmprojout_7_dataarray_data_V_ce0       => open,
      vmprojout_7_dataarray_data_V_we0       => VMPROJ_24_mem_A_wea(L6PHIB16),
      vmprojout_7_dataarray_data_V_address0  => VMPROJ_24_mem_AV_writeaddr(L6PHIB16),
      vmprojout_7_dataarray_data_V_d0        => VMPROJ_24_mem_AV_din(L6PHIB16)
  );

  MC_start <= '1' when ME_done = '1';

  ME_L3PHIB9 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => ME_done,
      bx_V          => PR_bx_out,
      bx_o_V        => ME_bx_out,
      bx_o_V_ap_vld => ME_bx_out_vld,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB9n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB9n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB9n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB9n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB9),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB9),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB9),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB9)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB9)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB9),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB9),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB9)
  );

  ME_L3PHIB10 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB10n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB10n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB10n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB10n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB10),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB10),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB10),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB10)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB10)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB10),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB10),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB10)
  );

  ME_L3PHIB11 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB11n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB11n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB11n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB11n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB11),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB11),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB11),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB11)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB11)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB11),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB11),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB11)
  );

  ME_L3PHIB12 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB12n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB12n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB12n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB12n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB12),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB12),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB12),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB12)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB12)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB12),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB12),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB12)
  );

  ME_L3PHIB13 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB13n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB13n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB13n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB13n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB13),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB13),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB13),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB13)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB13)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB13),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB13),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB13)
  );

  ME_L3PHIB14 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB14n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB14n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB14n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB14n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB14),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB14),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB14),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB14)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB14)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB14),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB14),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB14)
  );

  ME_L3PHIB15 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB15n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB15n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB15n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB15n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB15),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB15),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB15),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB15)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB15)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB15),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB15),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB15)
  );

  ME_L3PHIB16 : entity work.ME_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_16_mem_A_enb(L3PHIB16n1),
      inputStubData_dataarray_data_V_address0  => VMSME_16_mem_AV_readaddr(L3PHIB16n1),
      inputStubData_dataarray_data_V_q0        => VMSME_16_mem_AV_dout(L3PHIB16n1),
      inputStubData_nentries_0_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_16_mem_AAAV_dout_nent(L3PHIB16n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L3PHIB16),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L3PHIB16),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L3PHIB16),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB16)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L3PHIB16)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L3PHIB16),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L3PHIB16),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L3PHIB16)
  );

  ME_L4PHIB9 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB9n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB9n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB9n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB9n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB9),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB9),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB9),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB9)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB9)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB9),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB9),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB9)
  );

  ME_L4PHIB10 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB10n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB10n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB10n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB10n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB10),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB10),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB10),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB10)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB10)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB10),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB10),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB10)
  );

  ME_L4PHIB11 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB11n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB11n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB11n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB11n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB11),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB11),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB11),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB11)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB11)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB11),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB11),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB11)
  );

  ME_L4PHIB12 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB12n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB12n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB12n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB12n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB12),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB12),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB12),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB12)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB12)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB12),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB12),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB12)
  );

  ME_L4PHIB13 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB13n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB13n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB13n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB13n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB13),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB13),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB13),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB13)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB13)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB13),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB13),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB13)
  );

  ME_L4PHIB14 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB14n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB14n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB14n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB14n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB14),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB14),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB14),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB14)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB14)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB14),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB14),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB14)
  );

  ME_L4PHIB15 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB15n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB15n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB15n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB15n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB15),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB15),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB15),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB15)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB15)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB15),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB15),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB15)
  );

  ME_L4PHIB16 : entity work.ME_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L4PHIB16n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L4PHIB16n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L4PHIB16n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L4PHIB16n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L4PHIB16),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L4PHIB16),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L4PHIB16),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB16)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L4PHIB16)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L4PHIB16),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L4PHIB16),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L4PHIB16)
  );

  ME_L5PHIB9 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB9n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB9n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB9n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB9n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB9),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB9),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB9),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB9)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB9)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB9),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB9),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB9)
  );

  ME_L5PHIB10 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB10n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB10n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB10n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB10n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB10),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB10),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB10),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB10)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB10)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB10),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB10),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB10)
  );

  ME_L5PHIB11 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB11n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB11n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB11n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB11n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB11),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB11),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB11),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB11)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB11)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB11),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB11),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB11)
  );

  ME_L5PHIB12 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB12n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB12n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB12n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB12n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB12),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB12),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB12),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB12)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB12)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB12),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB12),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB12)
  );

  ME_L5PHIB13 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB13n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB13n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB13n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB13n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB13),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB13),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB13),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB13)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB13)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB13),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB13),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB13)
  );

  ME_L5PHIB14 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB14n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB14n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB14n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB14n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB14),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB14),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB14),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB14)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB14)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB14),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB14),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB14)
  );

  ME_L5PHIB15 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB15n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB15n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB15n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB15n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB15),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB15),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB15),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB15)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB15)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB15),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB15),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB15)
  );

  ME_L5PHIB16 : entity work.ME_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L5PHIB16n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L5PHIB16n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L5PHIB16n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L5PHIB16n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L5PHIB16),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L5PHIB16),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L5PHIB16),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB16)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L5PHIB16)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L5PHIB16),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L5PHIB16),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L5PHIB16)
  );

  ME_L6PHIB9 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB9n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB9n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB9n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB9n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB9),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB9),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB9),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB9)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB9)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB9),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB9),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB9)
  );

  ME_L6PHIB10 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB10n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB10n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB10n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB10n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB10),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB10),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB10),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB10)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB10)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB10),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB10),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB10)
  );

  ME_L6PHIB11 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB11n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB11n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB11n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB11n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB11),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB11),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB11),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB11)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB11)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB11),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB11),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB11)
  );

  ME_L6PHIB12 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB12n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB12n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB12n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB12n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB12),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB12),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB12),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB12)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB12)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB12),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB12),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB12)
  );

  ME_L6PHIB13 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB13n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB13n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB13n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB13n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB13),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB13),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB13),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB13)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB13)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB13),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB13),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB13)
  );

  ME_L6PHIB14 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB14n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB14n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB14n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB14n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB14),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB14),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB14),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB14)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB14)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB14),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB14),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB14)
  );

  ME_L6PHIB15 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB15n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB15n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB15n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB15n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB15),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB15),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB15),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB15)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB15)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB15),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB15),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB15)
  );

  ME_L6PHIB16 : entity work.ME_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => ME_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => PR_bx_out,
      inputStubData_dataarray_data_V_ce0       => VMSME_17_mem_A_enb(L6PHIB16n1),
      inputStubData_dataarray_data_V_address0  => VMSME_17_mem_AV_readaddr(L6PHIB16n1),
      inputStubData_dataarray_data_V_q0        => VMSME_17_mem_AV_dout(L6PHIB16n1),
      inputStubData_nentries_0_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(0),
      inputStubData_nentries_0_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(1),
      inputStubData_nentries_0_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(2),
      inputStubData_nentries_0_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(3),
      inputStubData_nentries_0_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(4),
      inputStubData_nentries_0_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(5),
      inputStubData_nentries_0_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(6),
      inputStubData_nentries_0_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(0)(7),
      inputStubData_nentries_1_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(0),
      inputStubData_nentries_1_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(1),
      inputStubData_nentries_1_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(2),
      inputStubData_nentries_1_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(3),
      inputStubData_nentries_1_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(4),
      inputStubData_nentries_1_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(5),
      inputStubData_nentries_1_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(6),
      inputStubData_nentries_1_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(1)(7),
      inputStubData_nentries_2_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(0),
      inputStubData_nentries_2_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(1),
      inputStubData_nentries_2_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(2),
      inputStubData_nentries_2_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(3),
      inputStubData_nentries_2_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(4),
      inputStubData_nentries_2_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(5),
      inputStubData_nentries_2_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(6),
      inputStubData_nentries_2_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(2)(7),
      inputStubData_nentries_3_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(0),
      inputStubData_nentries_3_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(1),
      inputStubData_nentries_3_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(2),
      inputStubData_nentries_3_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(3),
      inputStubData_nentries_3_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(4),
      inputStubData_nentries_3_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(5),
      inputStubData_nentries_3_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(6),
      inputStubData_nentries_3_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(3)(7),
      inputStubData_nentries_4_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(0),
      inputStubData_nentries_4_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(1),
      inputStubData_nentries_4_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(2),
      inputStubData_nentries_4_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(3),
      inputStubData_nentries_4_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(4),
      inputStubData_nentries_4_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(5),
      inputStubData_nentries_4_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(6),
      inputStubData_nentries_4_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(4)(7),
      inputStubData_nentries_5_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(0),
      inputStubData_nentries_5_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(1),
      inputStubData_nentries_5_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(2),
      inputStubData_nentries_5_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(3),
      inputStubData_nentries_5_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(4),
      inputStubData_nentries_5_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(5),
      inputStubData_nentries_5_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(6),
      inputStubData_nentries_5_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(5)(7),
      inputStubData_nentries_6_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(0),
      inputStubData_nentries_6_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(1),
      inputStubData_nentries_6_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(2),
      inputStubData_nentries_6_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(3),
      inputStubData_nentries_6_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(4),
      inputStubData_nentries_6_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(5),
      inputStubData_nentries_6_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(6),
      inputStubData_nentries_6_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(6)(7),
      inputStubData_nentries_7_V_0     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(0),
      inputStubData_nentries_7_V_1     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(1),
      inputStubData_nentries_7_V_2     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(2),
      inputStubData_nentries_7_V_3     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(3),
      inputStubData_nentries_7_V_4     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(4),
      inputStubData_nentries_7_V_5     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(5),
      inputStubData_nentries_7_V_6     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(6),
      inputStubData_nentries_7_V_7     => VMSME_17_mem_AAAV_dout_nent(L6PHIB16n1)(7)(7),
      inputProjectionData_dataarray_data_V_ce0       => VMPROJ_24_mem_A_enb(L6PHIB16),
      inputProjectionData_dataarray_data_V_address0  => VMPROJ_24_mem_AV_readaddr(L6PHIB16),
      inputProjectionData_dataarray_data_V_q0        => VMPROJ_24_mem_AV_dout(L6PHIB16),
      inputProjectionData_nentries_0_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB16)(0),
      inputProjectionData_nentries_1_V               => VMPROJ_24_mem_AAV_dout_nent(L6PHIB16)(1),
      outputCandidateMatch_dataarray_data_V_ce0       => open,
      outputCandidateMatch_dataarray_data_V_we0       => CM_14_mem_A_wea(L6PHIB16),
      outputCandidateMatch_dataarray_data_V_address0  => CM_14_mem_AV_writeaddr(L6PHIB16),
      outputCandidateMatch_dataarray_data_V_d0        => CM_14_mem_AV_din(L6PHIB16)
  );

  FT_start <= '1' when MC_done = '1';

  MC_L3PHIB : entity work.MC_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => MC_done,
      bx_V          => ME_bx_out,
      bx_o_V        => MC_bx_out,
      bx_o_V_ap_vld => MC_bx_out_vld,
      match_0_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB9),
      match_0_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB9),
      match_0_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB9),
      match_0_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB9)(0),
      match_0_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB9)(1),
      match_1_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB10),
      match_1_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB10),
      match_1_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB10),
      match_1_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB10)(0),
      match_1_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB10)(1),
      match_2_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB11),
      match_2_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB11),
      match_2_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB11),
      match_2_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB11)(0),
      match_2_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB11)(1),
      match_3_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB12),
      match_3_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB12),
      match_3_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB12),
      match_3_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB12)(0),
      match_3_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB12)(1),
      match_4_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB13),
      match_4_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB13),
      match_4_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB13),
      match_4_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB13)(0),
      match_4_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB13)(1),
      match_5_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB14),
      match_5_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB14),
      match_5_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB14),
      match_5_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB14)(0),
      match_5_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB14)(1),
      match_6_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB15),
      match_6_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB15),
      match_6_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB15),
      match_6_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB15)(0),
      match_6_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB15)(1),
      match_7_dataarray_data_V_ce0       => CM_14_mem_A_enb(L3PHIB16),
      match_7_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L3PHIB16),
      match_7_dataarray_data_V_q0        => CM_14_mem_AV_dout(L3PHIB16),
      match_7_nentries_0_V               => CM_14_mem_AAV_dout_nent(L3PHIB16)(0),
      match_7_nentries_1_V               => CM_14_mem_AAV_dout_nent(L3PHIB16)(1),
      allstub_dataarray_data_V_ce0       => AS_36_mem_A_enb(L3PHIBn1),
      allstub_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L3PHIBn1),
      allstub_dataarray_data_V_q0        => AS_36_mem_AV_dout(L3PHIBn1),
      allproj_dataarray_data_V_ce0       => AP_60_mem_A_enb(L3PHIB),
      allproj_dataarray_data_V_address0  => AP_60_mem_AV_readaddr(L3PHIB),
      allproj_dataarray_data_V_q0        => AP_60_mem_AV_dout(L3PHIB),
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_52_mem_A_wea(L1L2_L3PHIB),
      fullmatch_0_dataarray_data_V_address0  => FM_52_mem_AV_writeaddr(L1L2_L3PHIB),
      fullmatch_0_dataarray_data_V_d0        => FM_52_mem_AV_din(L1L2_L3PHIB)
  );

  MC_L4PHIB : entity work.MC_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => ME_bx_out,
      match_0_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB9),
      match_0_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB9),
      match_0_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB9),
      match_0_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB9)(0),
      match_0_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB9)(1),
      match_1_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB10),
      match_1_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB10),
      match_1_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB10),
      match_1_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB10)(0),
      match_1_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB10)(1),
      match_2_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB11),
      match_2_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB11),
      match_2_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB11),
      match_2_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB11)(0),
      match_2_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB11)(1),
      match_3_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB12),
      match_3_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB12),
      match_3_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB12),
      match_3_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB12)(0),
      match_3_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB12)(1),
      match_4_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB13),
      match_4_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB13),
      match_4_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB13),
      match_4_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB13)(0),
      match_4_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB13)(1),
      match_5_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB14),
      match_5_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB14),
      match_5_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB14),
      match_5_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB14)(0),
      match_5_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB14)(1),
      match_6_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB15),
      match_6_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB15),
      match_6_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB15),
      match_6_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB15)(0),
      match_6_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB15)(1),
      match_7_dataarray_data_V_ce0       => CM_14_mem_A_enb(L4PHIB16),
      match_7_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L4PHIB16),
      match_7_dataarray_data_V_q0        => CM_14_mem_AV_dout(L4PHIB16),
      match_7_nentries_0_V               => CM_14_mem_AAV_dout_nent(L4PHIB16)(0),
      match_7_nentries_1_V               => CM_14_mem_AAV_dout_nent(L4PHIB16)(1),
      allstub_dataarray_data_V_ce0       => AS_36_mem_A_enb(L4PHIBn1),
      allstub_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L4PHIBn1),
      allstub_dataarray_data_V_q0        => AS_36_mem_AV_dout(L4PHIBn1),
      allproj_dataarray_data_V_ce0       => AP_58_mem_A_enb(L4PHIB),
      allproj_dataarray_data_V_address0  => AP_58_mem_AV_readaddr(L4PHIB),
      allproj_dataarray_data_V_q0        => AP_58_mem_AV_dout(L4PHIB),
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_52_mem_A_wea(L1L2_L4PHIB),
      fullmatch_0_dataarray_data_V_address0  => FM_52_mem_AV_writeaddr(L1L2_L4PHIB),
      fullmatch_0_dataarray_data_V_d0        => FM_52_mem_AV_din(L1L2_L4PHIB)
  );

  MC_L5PHIB : entity work.MC_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => ME_bx_out,
      match_0_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB9),
      match_0_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB9),
      match_0_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB9),
      match_0_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB9)(0),
      match_0_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB9)(1),
      match_1_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB10),
      match_1_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB10),
      match_1_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB10),
      match_1_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB10)(0),
      match_1_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB10)(1),
      match_2_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB11),
      match_2_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB11),
      match_2_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB11),
      match_2_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB11)(0),
      match_2_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB11)(1),
      match_3_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB12),
      match_3_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB12),
      match_3_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB12),
      match_3_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB12)(0),
      match_3_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB12)(1),
      match_4_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB13),
      match_4_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB13),
      match_4_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB13),
      match_4_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB13)(0),
      match_4_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB13)(1),
      match_5_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB14),
      match_5_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB14),
      match_5_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB14),
      match_5_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB14)(0),
      match_5_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB14)(1),
      match_6_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB15),
      match_6_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB15),
      match_6_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB15),
      match_6_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB15)(0),
      match_6_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB15)(1),
      match_7_dataarray_data_V_ce0       => CM_14_mem_A_enb(L5PHIB16),
      match_7_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L5PHIB16),
      match_7_dataarray_data_V_q0        => CM_14_mem_AV_dout(L5PHIB16),
      match_7_nentries_0_V               => CM_14_mem_AAV_dout_nent(L5PHIB16)(0),
      match_7_nentries_1_V               => CM_14_mem_AAV_dout_nent(L5PHIB16)(1),
      allstub_dataarray_data_V_ce0       => AS_36_mem_A_enb(L5PHIBn1),
      allstub_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L5PHIBn1),
      allstub_dataarray_data_V_q0        => AS_36_mem_AV_dout(L5PHIBn1),
      allproj_dataarray_data_V_ce0       => AP_58_mem_A_enb(L5PHIB),
      allproj_dataarray_data_V_address0  => AP_58_mem_AV_readaddr(L5PHIB),
      allproj_dataarray_data_V_q0        => AP_58_mem_AV_dout(L5PHIB),
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_52_mem_A_wea(L1L2_L5PHIB),
      fullmatch_0_dataarray_data_V_address0  => FM_52_mem_AV_writeaddr(L1L2_L5PHIB),
      fullmatch_0_dataarray_data_V_d0        => FM_52_mem_AV_din(L1L2_L5PHIB)
  );

  MC_L6PHIB : entity work.MC_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => ME_bx_out,
      match_0_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB9),
      match_0_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB9),
      match_0_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB9),
      match_0_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB9)(0),
      match_0_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB9)(1),
      match_1_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB10),
      match_1_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB10),
      match_1_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB10),
      match_1_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB10)(0),
      match_1_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB10)(1),
      match_2_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB11),
      match_2_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB11),
      match_2_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB11),
      match_2_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB11)(0),
      match_2_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB11)(1),
      match_3_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB12),
      match_3_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB12),
      match_3_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB12),
      match_3_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB12)(0),
      match_3_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB12)(1),
      match_4_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB13),
      match_4_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB13),
      match_4_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB13),
      match_4_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB13)(0),
      match_4_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB13)(1),
      match_5_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB14),
      match_5_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB14),
      match_5_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB14),
      match_5_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB14)(0),
      match_5_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB14)(1),
      match_6_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB15),
      match_6_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB15),
      match_6_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB15),
      match_6_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB15)(0),
      match_6_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB15)(1),
      match_7_dataarray_data_V_ce0       => CM_14_mem_A_enb(L6PHIB16),
      match_7_dataarray_data_V_address0  => CM_14_mem_AV_readaddr(L6PHIB16),
      match_7_dataarray_data_V_q0        => CM_14_mem_AV_dout(L6PHIB16),
      match_7_nentries_0_V               => CM_14_mem_AAV_dout_nent(L6PHIB16)(0),
      match_7_nentries_1_V               => CM_14_mem_AAV_dout_nent(L6PHIB16)(1),
      allstub_dataarray_data_V_ce0       => AS_36_mem_A_enb(L6PHIBn1),
      allstub_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L6PHIBn1),
      allstub_dataarray_data_V_q0        => AS_36_mem_AV_dout(L6PHIBn1),
      allproj_dataarray_data_V_ce0       => AP_58_mem_A_enb(L6PHIB),
      allproj_dataarray_data_V_address0  => AP_58_mem_AV_readaddr(L6PHIB),
      allproj_dataarray_data_V_q0        => AP_58_mem_AV_dout(L6PHIB),
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_52_mem_A_wea(L1L2_L6PHIB),
      fullmatch_0_dataarray_data_V_address0  => FM_52_mem_AV_writeaddr(L1L2_L6PHIB),
      fullmatch_0_dataarray_data_V_d0        => FM_52_mem_AV_din(L1L2_L6PHIB)
  );

  FT_L1L2 : entity work.FT_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => FT_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => FT_done,
      bx_V          => MC_bx_out,
      bx_o_V        => FT_bx_out,
      bx_o_V_ap_vld => FT_bx_out_vld,
      trackletParameters_0_dataarray_data_V_ce0       => TPAR_70_mem_A_enb(L1L2F),
      trackletParameters_0_dataarray_data_V_address0  => TPAR_70_mem_AV_readaddr(L1L2F),
      trackletParameters_0_dataarray_data_V_q0        => TPAR_70_mem_AV_dout(L1L2F),
      barrelFullMatches_0_dataarray_data_V_ce0       => FM_52_mem_A_enb(L1L2_L3PHIB),
      barrelFullMatches_0_dataarray_data_V_address0  => FM_52_mem_AV_readaddr(L1L2_L3PHIB),
      barrelFullMatches_0_dataarray_data_V_q0        => FM_52_mem_AV_dout(L1L2_L3PHIB),
      barrelFullMatches_0_nentries_0_V               => FM_52_mem_AAV_dout_nent(L1L2_L3PHIB)(0),
      barrelFullMatches_0_nentries_1_V               => FM_52_mem_AAV_dout_nent(L1L2_L3PHIB)(1),
      barrelFullMatches_0_dataarray_data_V_ce1       => FM_52_mem_A_enb(L1L2_L3PHIB),
      barrelFullMatches_0_dataarray_data_V_address1  => FM_52_mem_AV_readaddr(L1L2_L3PHIB),
      barrelFullMatches_0_dataarray_data_V_q1        => FM_52_mem_AV_dout(L1L2_L3PHIB),
      barrelFullMatches_1_dataarray_data_V_ce0       => FM_52_mem_A_enb(L1L2_L4PHIB),
      barrelFullMatches_1_dataarray_data_V_address0  => FM_52_mem_AV_readaddr(L1L2_L4PHIB),
      barrelFullMatches_1_dataarray_data_V_q0        => FM_52_mem_AV_dout(L1L2_L4PHIB),
      barrelFullMatches_1_nentries_0_V               => FM_52_mem_AAV_dout_nent(L1L2_L4PHIB)(0),
      barrelFullMatches_1_nentries_1_V               => FM_52_mem_AAV_dout_nent(L1L2_L4PHIB)(1),
      barrelFullMatches_1_dataarray_data_V_ce1       => FM_52_mem_A_enb(L1L2_L4PHIB),
      barrelFullMatches_1_dataarray_data_V_address1  => FM_52_mem_AV_readaddr(L1L2_L4PHIB),
      barrelFullMatches_1_dataarray_data_V_q1        => FM_52_mem_AV_dout(L1L2_L4PHIB),
      barrelFullMatches_2_dataarray_data_V_ce0       => FM_52_mem_A_enb(L1L2_L5PHIB),
      barrelFullMatches_2_dataarray_data_V_address0  => FM_52_mem_AV_readaddr(L1L2_L5PHIB),
      barrelFullMatches_2_dataarray_data_V_q0        => FM_52_mem_AV_dout(L1L2_L5PHIB),
      barrelFullMatches_2_nentries_0_V               => FM_52_mem_AAV_dout_nent(L1L2_L5PHIB)(0),
      barrelFullMatches_2_nentries_1_V               => FM_52_mem_AAV_dout_nent(L1L2_L5PHIB)(1),
      barrelFullMatches_2_dataarray_data_V_ce1       => FM_52_mem_A_enb(L1L2_L5PHIB),
      barrelFullMatches_2_dataarray_data_V_address1  => FM_52_mem_AV_readaddr(L1L2_L5PHIB),
      barrelFullMatches_2_dataarray_data_V_q1        => FM_52_mem_AV_dout(L1L2_L5PHIB),
      barrelFullMatches_3_dataarray_data_V_ce0       => FM_52_mem_A_enb(L1L2_L6PHIB),
      barrelFullMatches_3_dataarray_data_V_address0  => FM_52_mem_AV_readaddr(L1L2_L6PHIB),
      barrelFullMatches_3_dataarray_data_V_q0        => FM_52_mem_AV_dout(L1L2_L6PHIB),
      barrelFullMatches_3_nentries_0_V               => FM_52_mem_AAV_dout_nent(L1L2_L6PHIB)(0),
      barrelFullMatches_3_nentries_1_V               => FM_52_mem_AAV_dout_nent(L1L2_L6PHIB)(1),
      barrelFullMatches_3_dataarray_data_V_ce1       => FM_52_mem_A_enb(L1L2_L6PHIB),
      barrelFullMatches_3_dataarray_data_V_address1  => FM_52_mem_AV_readaddr(L1L2_L6PHIB),
      barrelFullMatches_3_dataarray_data_V_q1        => FM_52_mem_AV_dout(L1L2_L6PHIB),
      trackWord_V_din       => TW_84_stream_AV_din(L1L2),
      trackWord_V_full_n    => TW_84_stream_A_full_neg(L1L2),
      trackWord_V_write     => TW_84_stream_A_write(L1L2),
      barrelStubWords_0_V_din       => BW_46_stream_AV_din(L1L2_L3),
      barrelStubWords_0_V_full_n    => BW_46_stream_A_full_neg(L1L2_L3),
      barrelStubWords_0_V_write     => BW_46_stream_A_write(L1L2_L3),
      barrelStubWords_1_V_din       => BW_46_stream_AV_din(L1L2_L4),
      barrelStubWords_1_V_full_n    => BW_46_stream_A_full_neg(L1L2_L4),
      barrelStubWords_1_V_write     => BW_46_stream_A_write(L1L2_L4),
      barrelStubWords_2_V_din       => BW_46_stream_AV_din(L1L2_L5),
      barrelStubWords_2_V_full_n    => BW_46_stream_A_full_neg(L1L2_L5),
      barrelStubWords_2_V_write     => BW_46_stream_A_write(L1L2_L5),
      barrelStubWords_3_V_din       => BW_46_stream_AV_din(L1L2_L6),
      barrelStubWords_3_V_full_n    => BW_46_stream_A_full_neg(L1L2_L6),
      barrelStubWords_3_V_write     => BW_46_stream_A_write(L1L2_L6)
  );



end rtl;
